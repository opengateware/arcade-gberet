//------------------------------------------------------------------------------
// SPDX-License-Identifier: GPL-3.0-or-later
// SPDX-FileType: SOURCE
// SPDX-FileCopyrightText: (c) 2013-2019 MiSTer-X
//------------------------------------------------------------------------------

`ifndef __HID_DEFINITION
`define __HID_DEFINITION

`define none  1'b0

`define COIN2 INP2[3]
`define COIN1 INP2[2]
`define P1ST  INP2[0]
`define P2ST  INP2[1]

`define P1UP  INP0[0]
`define P1DW  INP0[2]
`define P1LF  INP0[3]
`define P1RG  INP0[1]
`define P1TA  INP0[4]
`define P1TB  INP0[5]

`define P2UP  INP1[0]
`define P2DW  INP1[2]
`define P2LF  INP1[3]
`define P2RG  INP1[1]
`define P2TA  INP1[4]
`define P2TB  INP1[5]

`endif
